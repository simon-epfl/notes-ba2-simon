module updowncounter();


endmodule
